module hexfont
#( SIZE=64 )
( input wire [SIZE-1:0] in, output wire [(SIZE*2)-1:0] out );
	
	localparam DIGITS = SIZE / 4;
	
	genvar i;
	generate
		for (i = 0; i < DIGITS; i++) begin
			always_comb begin
				case(in[(i+1)*4-1:i*4])
					
					// +---+---+---+
					// |   | 6 |   |
					// +---+---+---+
					// | 1 |   | 5 |
					// +---+---+---+
					// |   | 0 |   |
					// +---+---+---+
					// | 2 |   | 4 |
					// +---+---+---+ +---+
					// |   | 3 |   | | 7 |
					// +---+---+---+ +---+
					
					4'h00: out[(i+1)*8-1:i*8] = 8'b01111110;
					4'h01: out[(i+1)*8-1:i*8] = 8'b00110000;
					4'h02: out[(i+1)*8-1:i*8] = 8'b01101101;
					4'h03: out[(i+1)*8-1:i*8] = 8'b01111001;
					4'h04: out[(i+1)*8-1:i*8] = 8'b00110011;
					4'h05: out[(i+1)*8-1:i*8] = 8'b01011011;
					4'h06: out[(i+1)*8-1:i*8] = 8'b01011111;
					4'h07: out[(i+1)*8-1:i*8] = 8'b01110000;
					4'h08: out[(i+1)*8-1:i*8] = 8'b01111111;
					4'h09: out[(i+1)*8-1:i*8] = 8'b01111011;
					4'h0a: out[(i+1)*8-1:i*8] = 8'b01110111;
					4'h0b: out[(i+1)*8-1:i*8] = 8'b00011111;
					4'h0c: out[(i+1)*8-1:i*8] = 8'b00001101;
					4'h0d: out[(i+1)*8-1:i*8] = 8'b00111101;
					4'h0e: out[(i+1)*8-1:i*8] = 8'b01001111;
					4'h0f: out[(i+1)*8-1:i*8] = 8'b01000111;
					default: out[(i+1)*8-1:i*8] = 8'b10000000; // DOT, never used.
				endcase
			end
		end
	endgenerate
endmodule

